primitive mux8_1 (Y, D0, D1, D2, D3, D4, D5, D6, D7, S2, S1, S0);
  output Y;
  input D0, D1, D2, D3, D4, D5, D6, D7, S2, S1, S0;

  table
    //D0 D1 D2 D3 D4 D5 D6 D7 S2 S1 S0 : Y
    ? ? ? ? ? ? ? ? x ? ? : x;
    ? ? ? ? ? ? ? ? ? x ? : x;
    ? ? ? ? ? ? ? ? ? ? x : x;

    //S=000 -> D0;
    0 ? ? ? ? ? ? ? 0 0 0 : 0;
    1 ? ? ? ? ? ? ? 0 0 0 : 1;

    //S=001 -> D1;
    ? 0 ? ? ? ? ? ? 0 0 1 : 0;
    ? 1 ? ? ? ? ? ? 0 0 1 : 1;

    //S=010 -> D2;
    ? ? 0 ? ? ? ? ? 0 1 0 : 0;
    ? ? 1 ? ? ? ? ? 0 1 0 : 1;

    //S=011 -> D3;
    ? ? ? 0 ? ? ? ? 0 1 1 : 0;
    ? ? ? 1 ? ? ? ? 0 1 1 : 1;

    //S=100 -> D4;
    ? ? ? ? 0 ? ? ? 1 0 0 : 0;
    ? ? ? ? 1 ? ? ? 1 0 0 : 1;

    //S=101 -> D5;
    ? ? ? ? ? 0 ? ? 1 0 1 : 0;
    ? ? ? ? ? 1 ? ? 1 0 1 : 1;

    //S=110 -> D6;
    ? ? ? ? ? ? 0 ? 1 1 0 : 0;
    ? ? ? ? ? ? 1 ? 1 1 0 : 1;

    //S=111 -> D7;
    ? ? ? ? ? ? ? 0 1 1 1 : 0;
    ? ? ? ? ? ? ? 1 1 1 1 : 1;

  endtable
endprimitive 

module mux8_1_TEST;
  reg [7:0] D;
  reg [2:0] S;
  wire Y;
  mux8_1 TF(Y, D[0], D[1], D[2], D[3], D[4], D[5], D[6], D[7], S[2], S[1], S[0]);

  initial begin
    $dumpfile("./out/wave.vcd");
    $dumpvars(0, mux8_1_TEST);

    $display(" D = 01011100");
    $display(" S[2:0] | Y |");
    $monitor(" %b    | %b |", S, Y);
    D=8'b01011100; S=3'b000; 

    #10 S=3'b001;
    #10 S=3'b010;
    #10 S=3'b011;
    #10 S=3'b100;
    #10 S=3'b101;
    #10 S=3'b110;
    #10 S=3'b111;

    #10 $finish;
  end
endmodule